library ieee;
use ieee.std_logic_1164.all;

entity lc_miniCPU is
    port(
        
    );
end entity lc_miniCPU;

architecture arch of lc_miniCPU is

end architecture arch;